/*
This file is part of verilog-buildingblocks,
by David R. Piegdon <dgit@piegdon.de>

verilog-buildingblocks is free software: you can redistribute it and/or modify
it under the terms of the GNU Lesser General Public License as published by
the Free Software Foundation, either version 3 of the License, or
(at your option) any later version.

verilog-buildingblocks is distributed in the hope that it will be useful,
but WITHOUT ANY WARRANTY; without even the implied warranty of
MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
GNU Lesser General Public License for more details.

You should have received a copy of the GNU Lesser General Public License
along with verilog-buildingblocks.  If not, see <https://www.gnu.org/licenses/>.
*/

`ifndef __vbb__lattice_ice40__pullup_input_v__
`define __vbb__lattice_ice40__pullup_input_v__

`default_nettype none

// Implementation of input with pullup.
module pullup_input(input pin, output wire value);
	SB_IO #(
		.PIN_TYPE(6'b0000_01),
		.PULLUP(1'b1),
	) sb_io (
		.PACKAGE_PIN(pin),
		.D_IN_0(value),
	);
endmodule

`endif // __vbb__lattice_ice40__pullup_input_v__
