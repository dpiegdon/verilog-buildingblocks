`default_nettype none

module fifo();

	parameter WIDTH 8;
	parameter DEPTH 16;

endmodule

